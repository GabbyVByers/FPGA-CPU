module KEYBOARD_PLACEHOLDER (
	output wire [15:0] KEY 
);

assign KEY = 16'd0;

endmodule

