module KEYBOARD_PLACEHOLDER (
	output wire [15:0] KEY 
);

// Placeholder
assign KEY = 16'd0;

endmodule


